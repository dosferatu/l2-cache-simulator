//**************************************************
// L2 Cache module
//
//**************************************************

module L2Cache(L1BusIn, L1BusOut, L1OperationBusIn, sharedBusIn, sharedBusOut, sharedOperationBusIn, sharedOperationOut, snoopBusIn, snoopBusOut, hit, miss, read, write);

/*************************************************************************************************************/
/*                                       This section establishes parameters                                 */
/*                                    and defines input/outputs for the module.                              */
/*                                        It also initializes variables for                                  */
/*                                                use by the module.                                         */
/*************************************************************************************************************/
  // Establish parameters that can be used for dynamic sizing of cache
  parameter addressSize     = 32;   // Instruction size used by architecture
  parameter byteSelectBits  = 6;    // Number of byte select bits according to line size
  parameter indexBits       = 14;   // Number of bits from the address used for indexing to a set in way
  parameter lineSize        = 512;  // Size of the line of data in a set and used for shared bus size
  parameter L1BusSize       = 256;  // Size of Bus to communicate with the L1
  parameter tagBits         = 12;   // Number of bits from the address used for tag for validating index
  parameter ways            = 8;    // Number of ways for set associativity
  parameter M               = 1;    //
  parameter E               = 2;    //
  parameter S               = 4;    //
  parameter I               = 8;    //  
  parameter display         = 0;    // Set display flag

  // Declare inputs and outputs
  input       [lineSize - 1:0]  sharedBusIn;
  output reg  [lineSize - 1:0]  sharedBusOut;
  input       [255:0]           L1BusIn;
  output reg  [255:0]           L1BusOut;
  input       [15:0]            L1OperationBusIn;
  input       [7:0]             sharedOperationBusIn;
  output reg  [7:0]             sharedOperationBusOut;
  input       [1:0]             snoopBusIn;
  output reg  [1:0]             snoopBusOut;

  output reg  [31:0]            hit;
  output reg  [31:0]            miss;
  output reg  [31:0]            read;
  output reg  [31:0]            write;

  // Establish regs/registers for use by the module
  reg [tagBits - 1:0]        addressTag;   // Current operation's tag from address
  reg [byteSelectBits - 1:0] byteSelect;   // Current byte select value
  reg [lineSize - 1:0]       cacheData;    // Data from the cache line being operated on
  reg [tagBits - 1:0]        cacheTag;     // Tag from the cache line being operated on
  reg                        hitFlag;      // Stores whether a hit has occurred or not
  reg                        readFlag;     // Stores whether we are doing a read or a write operation
  reg                        writeFlag;    // 
  reg [indexBits - 1:0]      index;        // Currently selected set
  reg [$clog2(ways) - 1:0]   selectedWay;  // Current operation's selected way according to LRU

  reg [ways - 1:0]           COMPARATOR_OUT;       
  reg [lineSize - 1:0]       MUX_OUT;

  initial begin
    // Initialize statistics
    hit   = 0;
    miss  = 0;
    read  = 0;
    write = 0;
  end
  
  
  
/*************************************************************************************************************/
/*                                       This section establishes the cache                                  */
/*                                    data structure as a two dimensional array                              */
/*                                        of structures with data mebers:                                    */
/*                                        cacheTag, cacheData, mesi, lru                                     */
/*************************************************************************************************************/
  
  // Cache line structure
  typedef struct {
    bit[tagBits - 1:0] cacheTag;
    bit[lineSize - 1:0] cacheData;
    bit[3:0] mesi;
    bit[$clog2(ways) - 1:0] lru;
  } line;  
  
  // Generate n ways using n structs x m sets
  line Storage[ways - 1:0][2**indexBits - 1:0];

  // Initialize the L2 cache storage to an empty and invalidated state
  initial begin
    automatic integer i,j;
    automatic integer sets = 2**indexBits;

    for (i = 0; i < ways; i = i + 1) begin
      for (j = 0; j < sets; j = j + 1) begin
        Storage[i][j].cacheTag = 0;
        Storage[i][j].cacheData = 0;
        Storage[i][j].mesi = I;
        Storage[i][j].lru = 0;
      end
    end
  end


/*************************************************************************************************************/
/*                                     This section establishes the comparator                               */
/*                                  and multiplexor that will be used to check for                           */
/*                                    hits and get the data from the data cache                              */
/*************************************************************************************************************/

  // Generate parameter "ways" amount of comparators
  genvar i;
  generate
    for (i = 0; i < ways; i = i + 1) begin
      Comparator #(tagBits) comparator(addressTag, Storage[i][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheTag, COMPARATOR_OUT[i]);
    end
  endgenerate

  // Instantiate our encoder for n ways
  Encoder #(ways) encoder(COMPARATOR_OUT, ENCODER_OUT);

  // Wire up the cache data lines to the bus for the multiplexor input
  //  This is set up to allow as much as many as 16 ways
  case (ways)
    8: Multiplexor #(ways)  multiplexor(.select(ENCODER_OUT),
        .in0(Storage[0][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in1(Storage[1][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in2(Storage[2][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in3(Storage[3][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in4(Storage[4][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in5(Storage[5][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in6(Storage[6][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in7(Storage[7][L1BusIn[byteSelectBits + indexBits - 1:0]].cacheData),
        .in8(0),
        .in9(0),
        .in10(0),
        .in11(0),
        .in12(0),
        .in13(0),
        .in14(0),
        .in15(0),
        .out(MUX_OUT));
  endcase


/*************************************************************************************************************/
/*                                     This section establishes has the                                      */
/*                                  operations that will occur dependent on                                  */
/*                                    the inputs and states of the cache                                     */
/*************************************************************************************************************/

  // Performs necessary tasks/functions depending on whether there is a read or right to the cache
  always@(L1BusIn, L1OperationBusIn, sharedBusIn, sharedOperationBusIn) begin

    // Command 0
    if (L1OperationBusIn == "DR") begin
      // Update the cache
      CheckForHit;
      ReadL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(L1OperationBusIn);
    end

    // Command 1
    else if (L1OperationBus == "DW") begin
      // Update the cache
      CheckForHit;
      WriteL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(L1OperationBus);
    end

    // Command 2
    else if (L1OperationBus == "IR") begin
      // Update the cache
      CheckForHit;
      ReadL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(L1OperationBus);
    end

    // Command 3
    else if (sharedOperationBus == "I") begin
      // Update the cache
      CheckForHit;
      ReadL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(sharedOperationBus);
    end

    // Command 4
    else if (sharedOperationBus == "R") begin
      // Update the cache
      CheckForHit;
      ReadL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(sharedOperationBus);
    end

    // Command 5
    else if (sharedOperationBus == "W") begin
      // Update the cache
      CheckForHit;
      ReadL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(sharedOperationBus);
    end

    // Command 6
    else if (sharedOperationBus == "M") begin
      // Update the cache
      CheckForHit;
      ReadL2Cache;
      UpdateLRU;
      if (display == 1)
        DisplayState(sharedOperationBus);
    end

    // Command 8
    else if (L1OperationBus == "CL")
      ClearL2;

    // Command 9
    else if (L1OperationBus == "PR") begin
      DisplayValid;
    end
  end



/*************************************************************************************************************/
/*                                    This section defines tasks that will                                   */
/*                                  will be used by the L2Cache module to perform                            */
/*                                      appropriate operations on the cache                                  */
/*                                        dependent upon the cache inputs                                    */
/*************************************************************************************************************/

  task DisplayState (input[15:0] operation); begin
    automatic integer i;
    automatic string mesiStatus;

    // Display all elements of the current operation
    $display("Command: %s", operation);
    $display("L1 Bus (Hex): %h", L1BusIn[addressSize - 1:0]);
    $display("Shared Bus (Hex): %h", sharedBus[addressSize - 1:0]);
    $display("Address Tag (Hex): %h",addressTag);
    $display("Byte Select (Decimal): %d",byteSelect);
    $display("Index (Decimal): %d", index);

    // Display whether a hit or a miss
    if (hitFlag) begin
      $display("Cache hit from way: %d", selectedWay);
    end

    else if (~hitFlag) begin
      $display("Cache miss from way: %d", selectedWay);
    end

    // Loop through each way and see what the MESI state is for each
    for (i = 0; i < ways; i = i + 1) begin
      case (Storage[i][index].mesi)
        M: mesiStatus = "M";
        E: mesiStatus = "E";
        S: mesiStatus = "S";
        I: mesiStatus = "I";
      endcase

      $display("Way: %d\tLRU Value: %d\tMESI status: %s", i, Storage[i][index].lru, mesiStatus);
    end

    $display("\n");
  end
  endtask

  /****************************************************************************/

  // Update the hit detection flag and set the selected way if necessary.
  task CheckForHit; begin
    input [lineSize - 1:0]  address;
    automatic integer i;
    
    // Disect address
    addressTag  <= address[addressSize - 1:byteSelectBits + indexBits];
    byteSelect  <= address[byteSelectBits - 1:0];
    index       <= address[byteSelectBits + indexBits - 1:byteSelectBits];
    
    // Initialize hitFlag
    hitFlag = 0;

    // Check for hit from comparator and the mesi bits of the ways
    for (i = 0; i < ways; i = i + 1) begin
      hitFlag = hitFlag | (COMPARATOR_OUT[i] & ~Storage[i][index].mesi[3]);
    end
    
    // Increment hits and misses
    if (hitFlag) begin
      hit         <= hit + 1;
      selectedWay <= ENCODER_OUT; 
    end
    else if (!hitFlag)
      miss = miss + 1;
  end
  endtask

/*********************************************************************/

  task WriteL2Cache; begin
    write = write + 1;

    if (hitFlag)
      Storage[selectedWay][index].cacheData <= "W";
    else if (!hitFlag) begin
      QueryLRU;
      case(Storage[selectedWay][index].mesi)
        M: begin
          WriteSharedBus;
          Storage[selectedWay][index].cachData = "W";
        end
        
        E: Storage[selectedWay][index].cachData = "W";

        S: Storage[selectedWay][index].cachData = "W";

        I: Storage[selectedWay][index].cachData = "W";
      end
    endcase
  end
  endtask
  
/****************************************************************************/

  task ReadL2Cache; begin
    read = read + 1;
    WriteL1;
  endtask

/***************************************************************/

  task ReadSharedBus; begin
    input [7:0]   operation;
    
    if(operation == "R") begin
      sharedOperationBusOut <= operation;
      sharedBusOut          <= address;
    end
    else if(operation == "M") begin
      sharedOperationBusOut <= operation;
      sharedBusOut          <= address;
    end
  endtask

/********************************************************************/

  task WriteSharedBus; begin
    input [lineSize - 1:0] address;
    reg   [lineSize - 1:0] newAddress;
    
    assign newAddress = address & 6'b000000;
    sharedBusOut          <= newAddress;
    sharedOperationBusOut <= "W";
  end
  endtask

/*********************************************************************/

  task WriteL1; begin
    if (sharedOperationBusIn == "I")
      L1BusOut <= sharedBusIn & 5'b00000;
    else if (L1OperationBusIn == "DR")
      L1BusOut <= "L1DR";
    else if (L1OperationBusIn == "DW")
      L1BusOut <= "L1DW";
    else
      L1BusOut <= "L1IR";
  end
  endtask

/*********************************************************************/

  task SendInvalidate; begin
    sharedBusOut        <= L1BusIn & 5'b00000;
    sharedOperationBus  <= "I";
  end
  endtask

/*********************************************************************/

  task InvalidateL2; begin
    input [lineSize - 1:0]  address;
    
    // Invalidate line
    Storage[selectedWay][address[byteSelectBits + indexBits - 1:byteSelectBits].mesi = "I";
    
    // Send L1 Bus address to invalidate     
    L1BusOut = address & 5'b00000;
  end
  endtask

/*********************************************************************/

  // Clear cache & reset all states
  task ClearL2; begin
    automatic integer i,j;
    automatic integer sets = 2**indexBits;

    for (i = 0; i < ways; i = i + 1) begin
      for (j = 0; j < sets; j = j + 1) begin
        Storage[i][j].mesi = I;
        Storage[i][j].lru = 0;
      end
    end
  end
  endtask

/*********************************************************************/

  // Print contents and state of each valid
  task DisplayValid; begin
    automatic integer i,j;
    automatic integer sets = 2**indexBits;
    
    for (i = 0; i < ways; i = i + 1) begin
      for (j = 0; j < sets; j = j + 1) begin
        if(Storage[i][j].mesi != I);
        $display("Way: %d \t Index: %h \t MESI: %b \t LRU: %d", i, j, Storage[i][j].mesi, Storage[i][j].lru);
      end
    end
    endtask

/*********************************************************************/

  // Loop through the set array at row[index]
  // Set the way to the least recently used column
  task QueryLRU; begin
    automatic integer LRUvalue = 0;
    automatic integer i;

    // Loop through each way to find which way is LRU
    // i is used to keep track of the current way during the loop
    for (i = 0;i < ways; i = i + 1) begin
      if (Storage[i][index].lru > LRUvalue) begin
        LRUvalue = Storage[i][index].lru;
        selectedWay = i;
      end
    end
  end
  endtask

/*********************************************************************/

  task UpdateLRU; begin
    automatic integer i;

    // Save the selected way's LRU value
    automatic reg[2:0] selectedLRU = Storage[selectedWay][index].lru;

    // Increment through each way at the index to check LRU values and update
    //  them accordingly
    for (i = 0; i < ways; i = i + 1) begin
      if (Storage[i][index].lru <= selectedLRU)
        Storage[i][index].lru = Storage[i][index].lru + 1;
    end

    // Finally set the selected way to the most recently used
    Storage[selectedWay][index].lru = 0;
    end
  endtask
  
/*********************************************************************/

  task PutSnoopResult; begin
    if (hitFlag) begin
      case(Storage[selectedWay][index].mesi)
        M: snoopBusout <= HITM;
        E: snoopBusOut <= HIT;
        S: snoopBusOut <= HIT;
        I: snoopBusOut <= MISS;
        default: snoopBusOut <= MISS;
    end
    else if(!hitFlag)
      snoopBusOut = MISS;
  end
  endtask
endmodule
