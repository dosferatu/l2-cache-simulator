module L2Cache(command, snoopBus, sharedBus);
  input command;
  output snoopBus, sharedBus;
end module
