library verilog;
use verilog.vl_types.all;
entity MESI_FSM_sv_unit is
end MESI_FSM_sv_unit;
