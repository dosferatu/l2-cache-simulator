//**************************************************
// Cache tag comparator:
// inputs: address tag, cache tag
// outputs: match
//**************************************************

module Comparator(
  addressTag[4:0],
  cacheTag[4:0],
  match
);

end module
