task convert;
  begin
    temp_out = (9/5) *( temp_in + 32);
  end
endtask
