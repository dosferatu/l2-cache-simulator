library verilog;
use verilog.vl_types.all;
entity FileIO_test is
end FileIO_test;
