library verilog;
use verilog.vl_types.all;
entity FSM_test is
end FSM_test;
