module ComparatorTestBench;
end module
