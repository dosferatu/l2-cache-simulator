library verilog;
use verilog.vl_types.all;
entity global_test_top is
end global_test_top;
