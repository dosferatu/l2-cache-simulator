library verilog;
use verilog.vl_types.all;
entity FSM_test_sv_unit is
end FSM_test_sv_unit;
